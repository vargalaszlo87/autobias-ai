* project: autobias-ai
* author: Varga Laszlo
* website: github.com/vargalaszlo87
*
* file: common emitter amplifier netlist
* version: 01
* last-updated:  2025.09.18

R1 N001 N005 {R1}
R2 N005 0 {R2}
RE N006 0 {RE}
RC N001 N002 {RC}
CE N006 0 {CE}
VCC N001 0 {VCC}
V1 N004 0 SINE(0 10m 1k)
CIN N005 N004 {CIN}
COUT out N002 {COUT}
RLOAD out 0 {RLOAD}

Q1 N002 N005 N006 0 QNPN
.model QNPN NPN (BF={HFE})

.options savecurrents
.temp 20
.fourier 1k V(out)
.param R1=10000 R2=2000 RC=1000 RE=0 CE=100u CIN=10u COUT=10u RLOAD=73 VCC=12 HFE=300
.control
op
tran 0.1m 20m 
wrdata output/tempFile.txt V(out) @RLOAD[i]
.endc
.end